-- Vhdl test bench created from schematic /home/karol/Desktop/UCISW/Projek1/test/pierwszy.sch - Fri Oct 24 02:30:46 2025
--
-- Notes: 
-- 1) This testbench template has been automatically generated using types
-- std_logic and std_logic_vector for the ports of the unit under test.
-- Xilinx recommends that these types always be used for the top-level
-- I/O of a design in order to guarantee that the testbench will bind
-- correctly to the timing (post-route) simulation model.
-- 2) To use this template as your testbench, change the filename to any
-- name of your choice with the extension .vhd, and use the "Source->Add"
-- menu in Project Navigator to import the testbench. Then
-- edit the user defined section below, adding code to generate the 
-- stimulus for your design.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY pierwszy_pierwszy_sch_tb IS
END pierwszy_pierwszy_sch_tb;
ARCHITECTURE behavioral OF pierwszy_pierwszy_sch_tb IS 

   COMPONENT pierwszy
   PORT( X	:	IN	STD_LOGIC_VECTOR (3 DOWNTO 0); 
          Y	:	OUT	STD_LOGIC_VECTOR (3 DOWNTO 0));
   END COMPONENT;

   SIGNAL X	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
   SIGNAL Y	:	STD_LOGIC_VECTOR (3 DOWNTO 0);

BEGIN

   UUT: pierwszy PORT MAP(
		X => X, 
		Y => Y
   );
	
		X <= "0000",
			"0001" after 200 ns,
			"1111" after 400 ns;

END;
